** Profile: "SCHEMATIC1-Bias"  [ C:\Documents and Settings\Javier\My Documents\EE10\PSpice 4\problem4-SCHEMATIC1-Bias.sim ] 

** Creating circuit file "problem4-SCHEMATIC1-Bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 500ms 0 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\problem4-SCHEMATIC1.net" 


.END
