APPLICATION CANCELED
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                           ;

		if (control = "0010" or control = "0011") then
				
			sel <= "10";

		end if;

		if (control = "1100" or control = "1110" or control = "1000" or control="1010") then
				
			sel <= "01";

		end if;


	end process;

end Behavioral;
