library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity dsadf is
    Port ( sdf : in std_logic_vector(15 downto 0));
end dsadf;

architecture Behavioral of dsadf is

begin


end Behavioral;
