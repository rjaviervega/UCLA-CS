** Profile: "SCHEMATIC1-Bias"  [ C:\DOCUMENTS AND SETTINGS\JAVIER\MY DOCUMENTS\EE10\PSpice 1\project 3-SCHEMATIC1-Bias.sim ] 

** Creating circuit file "project 3-SCHEMATIC1-Bias.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Program Files\OrcadLite\PSpice\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.PROBE V(*) I(*) W(*) D(*) NOISE(*) 
.INC ".\project 3-SCHEMATIC1.net" 


.END
