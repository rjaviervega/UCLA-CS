library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity shift is
    Port ( A : in std_logic_vector(15 downto 0);
           B : in std_logic_vector(3 downto 0);
           control : in std_logic_vector(3 downto 0);
           shift_result : out std_logic_vector(15 downto 0);
           shifted_out : out std_logic);
end shift;

architecture Behavioral of shift is

begin

	process (A, B, control) begin

	--- BEGIN sll, and sla

	-- Logical Shift
	if (control = "1100") then
		if B = "0000" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(14);
			shift_result(13) <= A(13);
			shift_result(12) <= A(12);
			shift_result(11) <= A(11);
			shift_result(10) <= A(10);
			shift_result(9) <= A(9);
			shift_result(8) <= A(8);
			shift_result(7) <= A(7);
			shift_result(6) <= A(6);
			shift_result(5) <= A(5);
			shift_result(4) <= A(4);
			shift_result(3) <= A(3);
			shift_result(2) <= A(2);
			shift_result(1) <= A(1);
			shift_result(0) <= A(0);
			shifted_out <= A(15);
		end if;
		if B = "0001" then
			shift_result(15) <= A(14);
			shift_result(14) <= A(13);
			shift_result(13) <= A(12);
			shift_result(12) <= A(11);
			shift_result(11) <= A(10);
			shift_result(10) <= A(9);
			shift_result(9) <= A(8);
			shift_result(8) <= A(7);
			shift_result(7) <= A(6);
			shift_result(6) <= A(5);
			shift_result(5) <= A(4);
			shift_result(4) <= A(3);
			shift_result(3) <= A(2);
			shift_result(2) <= A(1);
			shift_result(1) <= A(0);
			shift_result(0) <= '0';
			shifted_out <= A(15);
		end if;
		if B = "0010" then
			shift_result(15) <= A(13);
			shift_result(14) <= A(12);
			shift_result(13) <= A(11);
			shift_result(12) <= A(10);
			shift_result(11) <= A(9);
			shift_result(10) <= A(8);
			shift_result(9) <= A(7);
			shift_result(8) <= A(6);
			shift_result(7) <= A(5);
			shift_result(6) <= A(4);
			shift_result(5) <= A(3);
			shift_result(4) <= A(2);
			shift_result(3) <= A(1);
			shift_result(2) <= A(0);
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(14);
		end if;
		if B = "0011" then
			shift_result(15) <= A(12);
			shift_result(14) <= A(11);
			shift_result(13) <= A(10);
			shift_result(12) <= A(9);
			shift_result(11) <= A(8);
			shift_result(10) <= A(7);
			shift_result(9) <= A(6);
			shift_result(8) <= A(5);
			shift_result(7) <= A(4);
			shift_result(6) <= A(3);
			shift_result(5) <= A(2);
			shift_result(4) <= A(1);
			shift_result(3) <= A(0);
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(13);
		end if;
		if B = "0100" then
			shift_result(15) <= A(11);
			shift_result(14) <= A(10);
			shift_result(13) <= A(9);
			shift_result(12) <= A(8);
			shift_result(11) <= A(7);
			shift_result(10) <= A(6);
			shift_result(9) <= A(5);
			shift_result(8) <= A(4);
			shift_result(7) <= A(3);
			shift_result(6) <= A(2);
			shift_result(5) <= A(1);
			shift_result(4) <= A(0);
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(12);
		end if;
		if B = "0101" then
			shift_result(15) <= A(10);
			shift_result(14) <= A(9);
			shift_result(13) <= A(8);
			shift_result(12) <= A(7);
			shift_result(11) <= A(6);
			shift_result(10) <= A(5);
			shift_result(9) <= A(4);
			shift_result(8) <= A(3);
			shift_result(7) <= A(2);
			shift_result(6) <= A(1);
			shift_result(5) <= A(0);
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(11);
		end if;
		if B = "0110" then
			shift_result(15) <= A(9);
			shift_result(14) <= A(8);
			shift_result(13) <= A(7);
			shift_result(12) <= A(6);
			shift_result(11) <= A(5);
			shift_result(10) <= A(4);
			shift_result(9) <= A(3);
			shift_result(8) <= A(2);
			shift_result(7) <= A(1);
			shift_result(6) <= A(0);
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(10);
		end if;
		if B = "0111" then
			shift_result(15) <= A(8);
			shift_result(14) <= A(7);
			shift_result(13) <= A(6);
			shift_result(12) <= A(5);
			shift_result(11) <= A(4);
			shift_result(10) <= A(3);
			shift_result(9) <= A(2);
			shift_result(8) <= A(1);
			shift_result(7) <= A(0);
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(9);
		end if;
		if B = "1000" then
			shift_result(15) <= A(7);
			shift_result(14) <= A(6);
			shift_result(13) <= A(5);
			shift_result(12) <= A(4);
			shift_result(11) <= A(3);
			shift_result(10) <= A(2);
			shift_result(9) <= A(1);
			shift_result(8) <= A(0);
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(8);
		end if;
		if B = "1001" then
			shift_result(15) <= A(6);
			shift_result(14) <= A(5);
			shift_result(13) <= A(4);
			shift_result(12) <= A(3);
			shift_result(11) <= A(2);
			shift_result(10) <= A(1);
			shift_result(9) <= A(0);
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(7);
		end if;
		if B = "1010" then
			shift_result(15) <= A(5);
			shift_result(14) <= A(4);
			shift_result(13) <= A(3);
			shift_result(12) <= A(2);
			shift_result(11) <= A(1);
			shift_result(10) <= A(0);
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(6);
		end if;
		if B = "1011" then
			shift_result(15) <= A(4);
			shift_result(14) <= A(3);
			shift_result(13) <= A(2);
			shift_result(12) <= A(1);
			shift_result(11) <= A(0);
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(5);
		end if;
		if B = "1100" then
			shift_result(15) <= A(3);
			shift_result(14) <= A(2);
			shift_result(13) <= A(1);
			shift_result(12) <= A(0);
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(4);
		end if;
		if B = "1101" then
			shift_result(15) <= A(2);
			shift_result(14) <= A(1);
			shift_result(13) <= A(0);
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(3);
		end if;
		if B = "1110" then
			shift_result(15) <= A(1);
			shift_result(14) <= A(0);
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(2);
		end if;
		if B = "1111" then
			shift_result(15) <= A(0);
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(1);
		end if;
	end if;

	---  END sll, and sla

		
	--- BEGIN srl
	if control = "1110" then
		if B = "0000" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(14);
			shift_result(13) <= A(13);
			shift_result(12) <= A(12);
			shift_result(11) <= A(11);
			shift_result(10) <= A(10);
			shift_result(9) <= A(9);
			shift_result(8) <= A(8);
			shift_result(7) <= A(7);
			shift_result(6) <= A(6);
			shift_result(5) <= A(5);
			shift_result(4) <= A(4);
			shift_result(3) <= A(3);
			shift_result(2) <= A(2);
			shift_result(1) <= A(1);
			shift_result(0) <= A(0);
			shifted_out <= A(0);
		end if;
		if B = "0001" then
			shift_result(15) <= '0';
			shift_result(14) <= A(15);
			shift_result(13) <= A(14);
			shift_result(12) <= A(13);
			shift_result(11) <= A(12);
			shift_result(10) <= A(11);
			shift_result(9) <= A(10);
			shift_result(8) <= A(9);
			shift_result(7) <= A(8);
			shift_result(6) <= A(7);
			shift_result(5) <= A(6);
			shift_result(4) <= A(5);
			shift_result(3) <= A(4);
			shift_result(2) <= A(3);
			shift_result(1) <= A(2);
			shift_result(0) <= A(1);
			shifted_out <= A(0);
		end if;
		if B = "0010" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= A(15);
			shift_result(12) <= A(14);
			shift_result(11) <= A(13);
			shift_result(10) <= A(12);
			shift_result(9) <= A(11);
			shift_result(8) <= A(10);
			shift_result(7) <= A(9);
			shift_result(6) <= A(8);
			shift_result(5) <= A(7);
			shift_result(4) <= A(6);
			shift_result(3) <= A(5);
			shift_result(2) <= A(4);
			shift_result(1) <= A(3);
			shift_result(0) <= A(2);
			shifted_out <= A(1);
		end if;
		if B = "0011" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= A(15);
			shift_result(11) <= A(14);
			shift_result(10) <= A(13);
			shift_result(9) <= A(12);
			shift_result(8) <= A(11);
			shift_result(7) <= A(10);
			shift_result(6) <= A(9);
			shift_result(5) <= A(8);
			shift_result(4) <= A(7);
			shift_result(3) <= A(6);
			shift_result(2) <= A(5);
			shift_result(1) <= A(4);
			shift_result(0) <= A(3);
			shifted_out <= A(2);
		end if;
		if B = "0100" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= A(15);
			shift_result(10) <= A(14);
			shift_result(9) <= A(13);
			shift_result(8) <= A(12);
			shift_result(7) <= A(11);
			shift_result(6) <= A(10);
			shift_result(5) <= A(9);
			shift_result(4) <= A(8);
			shift_result(3) <= A(7);
			shift_result(2) <= A(6);
			shift_result(1) <= A(5);
			shift_result(0) <= A(4);
			shifted_out <= A(3);
		end if;
		if B = "0101" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= A(15);
			shift_result(9) <= A(14);
			shift_result(8) <= A(13);
			shift_result(7) <= A(12);
			shift_result(6) <= A(11);
			shift_result(5) <= A(10);
			shift_result(4) <= A(9);
			shift_result(3) <= A(8);
			shift_result(2) <= A(7);
			shift_result(1) <= A(6);
			shift_result(0) <= A(5);
			shifted_out <= A(4);
		end if;
		if B = "0110" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= A(15);
			shift_result(8) <= A(14);
			shift_result(7) <= A(13);
			shift_result(6) <= A(12);
			shift_result(5) <= A(11);
			shift_result(4) <= A(10);
			shift_result(3) <= A(9);
			shift_result(2) <= A(8);
			shift_result(1) <= A(7);
			shift_result(0) <= A(6);
			shifted_out <= A(5);
		end if;
		if B = "0111" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= A(15);
			shift_result(7) <= A(14);
			shift_result(6) <= A(13);
			shift_result(5) <= A(12);
			shift_result(4) <= A(11);
			shift_result(3) <= A(10);
			shift_result(2) <= A(9);
			shift_result(1) <= A(8);
			shift_result(0) <= A(7);
			shifted_out <= A(6);
		end if;
		if B = "1000" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= A(15);
			shift_result(6) <= A(14);
			shift_result(5) <= A(13);
			shift_result(4) <= A(12);
			shift_result(3) <= A(11);
			shift_result(2) <= A(10);
			shift_result(1) <= A(9);
			shift_result(0) <= A(8);
			shifted_out <= A(7);
		end if;
		if B = "1001" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= A(15);
			shift_result(5) <= A(14);
			shift_result(4) <= A(13);
			shift_result(3) <= A(12);
			shift_result(2) <= A(11);
			shift_result(1) <= A(10);
			shift_result(0) <= A(9);
			shifted_out <= A(8);
		end if;
		if B = "1010" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= A(15);
			shift_result(4) <= A(14);
			shift_result(3) <= A(13);
			shift_result(2) <= A(12);
			shift_result(1) <= A(11);
			shift_result(0) <= A(10);
			shifted_out <= A(9);
		end if;
		if B = "1011" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= A(15);
			shift_result(3) <= A(14);
			shift_result(2) <= A(13);
			shift_result(1) <= A(12);
			shift_result(0) <= A(11);
			shifted_out <= A(10);
		end if;
		if B = "1100" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= A(15);
			shift_result(2) <= A(14);
			shift_result(1) <= A(13);
			shift_result(0) <= A(12);
			shifted_out <= A(11);
		end if;
		if B = "1101" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= A(15);
			shift_result(1) <= A(14);
			shift_result(0) <= A(13);
			shifted_out <= A(12);
		end if;
		if B = "1110" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= A(15);
			shift_result(0) <= A(14);
			shifted_out <= A(13);
		end if;
		if B = "1111" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= A(15);
			shifted_out <= A(14);
		end if;
	end if;

	-- END srl

	-- BEGIN sla

	if control = "1010" then
		if B = "0000" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(14);
			shift_result(13) <= A(13);
			shift_result(12) <= A(12);
			shift_result(11) <= A(11);
			shift_result(10) <= A(10);
			shift_result(9) <= A(9);
			shift_result(8) <= A(8);
			shift_result(7) <= A(7);
			shift_result(6) <= A(6);
			shift_result(5) <= A(5);
			shift_result(4) <= A(4);
			shift_result(3) <= A(3);
			shift_result(2) <= A(2);
			shift_result(1) <= A(1);
			shift_result(0) <= A(0);
			shifted_out <= A(0);
		end if;
		if B = "0001" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(14);
			shift_result(12) <= A(13);
			shift_result(11) <= A(12);
			shift_result(10) <= A(11);
			shift_result(9) <= A(10);
			shift_result(8) <= A(9);
			shift_result(7) <= A(8);
			shift_result(6) <= A(7);
			shift_result(5) <= A(6);
			shift_result(4) <= A(5);
			shift_result(3) <= A(4);
			shift_result(2) <= A(3);
			shift_result(1) <= A(2);
			shift_result(0) <= A(1);
			shifted_out <= A(0);
		end if;
		if B = "0010" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(14);
			shift_result(11) <= A(13);
			shift_result(10) <= A(12);
			shift_result(9) <= A(11);
			shift_result(8) <= A(10);
			shift_result(7) <= A(9);
			shift_result(6) <= A(8);
			shift_result(5) <= A(7);
			shift_result(4) <= A(6);
			shift_result(3) <= A(5);
			shift_result(2) <= A(4);
			shift_result(1) <= A(3);
			shift_result(0) <= A(2);
			shifted_out <= A(1);
		end if;
		if B = "0011" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(14);
			shift_result(10) <= A(13);
			shift_result(9) <= A(12);
			shift_result(8) <= A(11);
			shift_result(7) <= A(10);
			shift_result(6) <= A(9);
			shift_result(5) <= A(8);
			shift_result(4) <= A(7);
			shift_result(3) <= A(6);
			shift_result(2) <= A(5);
			shift_result(1) <= A(4);
			shift_result(0) <= A(3);
			shifted_out <= A(2);
		end if;
		if B = "0100" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(14);
			shift_result(9) <= A(13);
			shift_result(8) <= A(12);
			shift_result(7) <= A(11);
			shift_result(6) <= A(10);
			shift_result(5) <= A(9);
			shift_result(4) <= A(8);
			shift_result(3) <= A(7);
			shift_result(2) <= A(6);
			shift_result(1) <= A(5);
			shift_result(0) <= A(4);
			shifted_out <= A(3);
		end if;
		if B = "0101" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(14);
			shift_result(8) <= A(13);
			shift_result(7) <= A(12);
			shift_result(6) <= A(11);
			shift_result(5) <= A(10);
			shift_result(4) <= A(9);
			shift_result(3) <= A(8);
			shift_result(2) <= A(7);
			shift_result(1) <= A(6);
			shift_result(0) <= A(5);
			shifted_out <= A(4);
		end if;
		if B = "0110" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(14);
			shift_result(7) <= A(13);
			shift_result(6) <= A(12);
			shift_result(5) <= A(11);
			shift_result(4) <= A(10);
			shift_result(3) <= A(9);
			shift_result(2) <= A(8);
			shift_result(1) <= A(7);
			shift_result(0) <= A(6);
			shifted_out <= A(5);
		end if;
		if B = "0111" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(14);
			shift_result(6) <= A(13);
			shift_result(5) <= A(12);
			shift_result(4) <= A(11);
			shift_result(3) <= A(10);
			shift_result(2) <= A(9);
			shift_result(1) <= A(8);
			shift_result(0) <= A(7);
			shifted_out <= A(6);
		end if;
		if B = "1000" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(14);
			shift_result(5) <= A(13);
			shift_result(4) <= A(12);
			shift_result(3) <= A(11);
			shift_result(2) <= A(10);
			shift_result(1) <= A(9);
			shift_result(0) <= A(8);
			shifted_out <= A(7);
		end if;
		if B = "1001" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(14);
			shift_result(4) <= A(13);
			shift_result(3) <= A(12);
			shift_result(2) <= A(11);
			shift_result(1) <= A(10);
			shift_result(0) <= A(9);
			shifted_out <= A(8);
		end if;
		if B = "1010" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(15);
			shift_result(4) <= A(14);
			shift_result(3) <= A(13);
			shift_result(2) <= A(12);
			shift_result(1) <= A(11);
			shift_result(0) <= A(10);
			shifted_out <= A(9);
		end if;
		if B = "1011" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(15);
			shift_result(4) <= A(15);
			shift_result(3) <= A(14);
			shift_result(2) <= A(13);
			shift_result(1) <= A(12);
			shift_result(0) <= A(11);
			shifted_out <= A(10);
		end if;
		if B = "1100" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(15);
			shift_result(4) <= A(15);
			shift_result(3) <= A(15);
			shift_result(2) <= A(14);
			shift_result(1) <= A(13);
			shift_result(0) <= A(12);
			shifted_out <= A(11);
		end if;
		if B = "1101" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(15);
			shift_result(4) <= A(15);
			shift_result(3) <= A(15);
			shift_result(2) <= A(15);
			shift_result(1) <= A(14);
			shift_result(0) <= A(13);
			shifted_out <= A(12);
		end if;
		if B = "1110" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(15);
			shift_result(4) <= A(15);
			shift_result(3) <= A(15);
			shift_result(2) <= A(15);
			shift_result(1) <= A(15);
			shift_result(0) <= A(14);
			shifted_out <= A(13);
		end if;
		if B = "1111" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(15);
			shift_result(4) <= A(15);
			shift_result(3) <= A(15);
			shift_result(2) <= A(15);
			shift_result(1) <= A(15);
			shift_result(0) <= A(15);
			shifted_out <= A(14);
		end if;
	end if;



	-- Arithm Shift
	if (control = "1000") then
		if B = "0000" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(14);
			shift_result(13) <= A(13);
			shift_result(12) <= A(12);
			shift_result(11) <= A(11);
			shift_result(10) <= A(10);
			shift_result(9) <= A(9);
			shift_result(8) <= A(8);
			shift_result(7) <= A(7);
			shift_result(6) <= A(6);
			shift_result(5) <= A(5);
			shift_result(4) <= A(4);
			shift_result(3) <= A(3);
			shift_result(2) <= A(2);
			shift_result(1) <= A(1);
			shift_result(0) <= A(0);
			shifted_out <= A(15);
		end if;
		if B = "0001" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(13);
			shift_result(13) <= A(12);
			shift_result(12) <= A(11);
			shift_result(11) <= A(10);
			shift_result(10) <= A(9);
			shift_result(9) <= A(8);
			shift_result(8) <= A(7);
			shift_result(7) <= A(6);
			shift_result(6) <= A(5);
			shift_result(5) <= A(4);
			shift_result(4) <= A(3);
			shift_result(3) <= A(2);
			shift_result(2) <= A(1);
			shift_result(1) <= A(0);
			shift_result(0) <= '0';
			shifted_out <= A(15);
		end if;
		if B = "0010" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(12);
			shift_result(13) <= A(11);
			shift_result(12) <= A(10);
			shift_result(11) <= A(9);
			shift_result(10) <= A(8);
			shift_result(9) <= A(7);
			shift_result(8) <= A(6);
			shift_result(7) <= A(5);
			shift_result(6) <= A(4);
			shift_result(5) <= A(3);
			shift_result(4) <= A(2);
			shift_result(3) <= A(1);
			shift_result(2) <= A(0);
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(14);
		end if;
		if B = "0011" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(11);
			shift_result(13) <= A(10);
			shift_result(12) <= A(9);
			shift_result(11) <= A(8);
			shift_result(10) <= A(7);
			shift_result(9) <= A(6);
			shift_result(8) <= A(5);
			shift_result(7) <= A(4);
			shift_result(6) <= A(3);
			shift_result(5) <= A(2);
			shift_result(4) <= A(1);
			shift_result(3) <= A(0);
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(13);
		end if;
		if B = "0100" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(10);
			shift_result(13) <= A(9);
			shift_result(12) <= A(8);
			shift_result(11) <= A(7);
			shift_result(10) <= A(6);
			shift_result(9) <= A(5);
			shift_result(8) <= A(4);
			shift_result(7) <= A(3);
			shift_result(6) <= A(2);
			shift_result(5) <= A(1);
			shift_result(4) <= A(0);
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(12);
		end if;
		if B = "0101" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(9);
			shift_result(13) <= A(8);
			shift_result(12) <= A(7);
			shift_result(11) <= A(6);
			shift_result(10) <= A(5);
			shift_result(9) <= A(4);
			shift_result(8) <= A(3);
			shift_result(7) <= A(2);
			shift_result(6) <= A(1);
			shift_result(5) <= A(0);
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(11);
		end if;
		if B = "0110" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(8);
			shift_result(13) <= A(7);
			shift_result(12) <= A(6);
			shift_result(11) <= A(5);
			shift_result(10) <= A(4);
			shift_result(9) <= A(3);
			shift_result(8) <= A(2);
			shift_result(7) <= A(1);
			shift_result(6) <= A(0);
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(10);
		end if;
		if B = "0111" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(7);
			shift_result(13) <= A(6);
			shift_result(12) <= A(5);
			shift_result(11) <= A(4);
			shift_result(10) <= A(3);
			shift_result(9) <= A(2);
			shift_result(8) <= A(1);
			shift_result(7) <= A(0);
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(9);
		end if;
		if B = "1000" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(6);
			shift_result(13) <= A(5);
			shift_result(12) <= A(4);
			shift_result(11) <= A(3);
			shift_result(10) <= A(2);
			shift_result(9) <= A(1);
			shift_result(8) <= A(0);
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(8);
		end if;
		if B = "1001" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(5);
			shift_result(13) <= A(4);
			shift_result(12) <= A(3);
			shift_result(11) <= A(2);
			shift_result(10) <= A(1);
			shift_result(9) <= A(0);
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(7);
		end if;
		if B = "1010" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(4);
			shift_result(13) <= A(3);
			shift_result(12) <= A(2);
			shift_result(11) <= A(1);
			shift_result(10) <= A(0);
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(6);
		end if;
		if B = "1011" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(3);
			shift_result(13) <= A(2);
			shift_result(12) <= A(1);
			shift_result(11) <= A(0);
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(5);
		end if;
		if B = "1100" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(2);
			shift_result(13) <= A(1);
			shift_result(12) <= A(0);
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(4);
		end if;
		if B = "1101" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(1);
			shift_result(13) <= A(0);
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(3);
		end if;
		if B = "1110" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(0);
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(2);
		end if;
		if B = "1111" then
			shift_result(15) <= A(15);
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= '0';
			shifted_out <= A(1);
		end if;
	end if;

	---  END sll, and sla

		
	--- BEGIN srl
	if control = "1110" then
		if B = "0000" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(14);
			shift_result(13) <= A(13);
			shift_result(12) <= A(12);
			shift_result(11) <= A(11);
			shift_result(10) <= A(10);
			shift_result(9) <= A(9);
			shift_result(8) <= A(8);
			shift_result(7) <= A(7);
			shift_result(6) <= A(6);
			shift_result(5) <= A(5);
			shift_result(4) <= A(4);
			shift_result(3) <= A(3);
			shift_result(2) <= A(2);
			shift_result(1) <= A(1);
			shift_result(0) <= A(0);
			shifted_out <= A(0);
		end if;
		if B = "0001" then
			shift_result(15) <= '0';
			shift_result(14) <= A(15);
			shift_result(13) <= A(14);
			shift_result(12) <= A(13);
			shift_result(11) <= A(12);
			shift_result(10) <= A(11);
			shift_result(9) <= A(10);
			shift_result(8) <= A(9);
			shift_result(7) <= A(8);
			shift_result(6) <= A(7);
			shift_result(5) <= A(6);
			shift_result(4) <= A(5);
			shift_result(3) <= A(4);
			shift_result(2) <= A(3);
			shift_result(1) <= A(2);
			shift_result(0) <= A(1);
			shifted_out <= A(0);
		end if;
		if B = "0010" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= A(15);
			shift_result(12) <= A(14);
			shift_result(11) <= A(13);
			shift_result(10) <= A(12);
			shift_result(9) <= A(11);
			shift_result(8) <= A(10);
			shift_result(7) <= A(9);
			shift_result(6) <= A(8);
			shift_result(5) <= A(7);
			shift_result(4) <= A(6);
			shift_result(3) <= A(5);
			shift_result(2) <= A(4);
			shift_result(1) <= A(3);
			shift_result(0) <= A(2);
			shifted_out <= A(1);
		end if;
		if B = "0011" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= A(15);
			shift_result(11) <= A(14);
			shift_result(10) <= A(13);
			shift_result(9) <= A(12);
			shift_result(8) <= A(11);
			shift_result(7) <= A(10);
			shift_result(6) <= A(9);
			shift_result(5) <= A(8);
			shift_result(4) <= A(7);
			shift_result(3) <= A(6);
			shift_result(2) <= A(5);
			shift_result(1) <= A(4);
			shift_result(0) <= A(3);
			shifted_out <= A(2);
		end if;
		if B = "0100" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= A(15);
			shift_result(10) <= A(14);
			shift_result(9) <= A(13);
			shift_result(8) <= A(12);
			shift_result(7) <= A(11);
			shift_result(6) <= A(10);
			shift_result(5) <= A(9);
			shift_result(4) <= A(8);
			shift_result(3) <= A(7);
			shift_result(2) <= A(6);
			shift_result(1) <= A(5);
			shift_result(0) <= A(4);
			shifted_out <= A(3);
		end if;
		if B = "0101" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= A(15);
			shift_result(9) <= A(14);
			shift_result(8) <= A(13);
			shift_result(7) <= A(12);
			shift_result(6) <= A(11);
			shift_result(5) <= A(10);
			shift_result(4) <= A(9);
			shift_result(3) <= A(8);
			shift_result(2) <= A(7);
			shift_result(1) <= A(6);
			shift_result(0) <= A(5);
			shifted_out <= A(4);
		end if;
		if B = "0110" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= A(15);
			shift_result(8) <= A(14);
			shift_result(7) <= A(13);
			shift_result(6) <= A(12);
			shift_result(5) <= A(11);
			shift_result(4) <= A(10);
			shift_result(3) <= A(9);
			shift_result(2) <= A(8);
			shift_result(1) <= A(7);
			shift_result(0) <= A(6);
			shifted_out <= A(5);
		end if;
		if B = "0111" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= A(15);
			shift_result(7) <= A(14);
			shift_result(6) <= A(13);
			shift_result(5) <= A(12);
			shift_result(4) <= A(11);
			shift_result(3) <= A(10);
			shift_result(2) <= A(9);
			shift_result(1) <= A(8);
			shift_result(0) <= A(7);
			shifted_out <= A(6);
		end if;
		if B = "1000" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= A(15);
			shift_result(6) <= A(14);
			shift_result(5) <= A(13);
			shift_result(4) <= A(12);
			shift_result(3) <= A(11);
			shift_result(2) <= A(10);
			shift_result(1) <= A(9);
			shift_result(0) <= A(8);
			shifted_out <= A(7);
		end if;
		if B = "1001" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= A(15);
			shift_result(5) <= A(14);
			shift_result(4) <= A(13);
			shift_result(3) <= A(12);
			shift_result(2) <= A(11);
			shift_result(1) <= A(10);
			shift_result(0) <= A(9);
			shifted_out <= A(8);
		end if;
		if B = "1010" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= A(15);
			shift_result(4) <= A(14);
			shift_result(3) <= A(13);
			shift_result(2) <= A(12);
			shift_result(1) <= A(11);
			shift_result(0) <= A(10);
			shifted_out <= A(9);
		end if;
		if B = "1011" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= A(15);
			shift_result(3) <= A(14);
			shift_result(2) <= A(13);
			shift_result(1) <= A(12);
			shift_result(0) <= A(11);
			shifted_out <= A(10);
		end if;
		if B = "1100" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= A(15);
			shift_result(2) <= A(14);
			shift_result(1) <= A(13);
			shift_result(0) <= A(12);
			shifted_out <= A(11);
		end if;
		if B = "1101" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= A(15);
			shift_result(1) <= A(14);
			shift_result(0) <= A(13);
			shifted_out <= A(12);
		end if;
		if B = "1110" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= A(15);
			shift_result(0) <= A(14);
			shifted_out <= A(13);
		end if;
		if B = "1111" then
			shift_result(15) <= '0';
			shift_result(14) <= '0';
			shift_result(13) <= '0';
			shift_result(12) <= '0';
			shift_result(11) <= '0';
			shift_result(10) <= '0';
			shift_result(9) <= '0';
			shift_result(8) <= '0';
			shift_result(7) <= '0';
			shift_result(6) <= '0';
			shift_result(5) <= '0';
			shift_result(4) <= '0';
			shift_result(3) <= '0';
			shift_result(2) <= '0';
			shift_result(1) <= '0';
			shift_result(0) <= A(15);
			shifted_out <= A(14);
		end if;
	end if;

	-- END srl

	-- BEGIN sla

	if control = "1010" then
		if B = "0000" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(14);
			shift_result(13) <= A(13);
			shift_result(12) <= A(12);
			shift_result(11) <= A(11);
			shift_result(10) <= A(10);
			shift_result(9) <= A(9);
			shift_result(8) <= A(8);
			shift_result(7) <= A(7);
			shift_result(6) <= A(6);
			shift_result(5) <= A(5);
			shift_result(4) <= A(4);
			shift_result(3) <= A(3);
			shift_result(2) <= A(2);
			shift_result(1) <= A(1);
			shift_result(0) <= A(0);
			shifted_out <= A(0);
		end if;
		if B = "0001" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(14);
			shift_result(12) <= A(13);
			shift_result(11) <= A(12);
			shift_result(10) <= A(11);
			shift_result(9) <= A(10);
			shift_result(8) <= A(9);
			shift_result(7) <= A(8);
			shift_result(6) <= A(7);
			shift_result(5) <= A(6);
			shift_result(4) <= A(5);
			shift_result(3) <= A(4);
			shift_result(2) <= A(3);
			shift_result(1) <= A(2);
			shift_result(0) <= A(1);
			shifted_out <= A(0);
		end if;
		if B = "0010" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(14);
			shift_result(11) <= A(13);
			shift_result(10) <= A(12);
			shift_result(9) <= A(11);
			shift_result(8) <= A(10);
			shift_result(7) <= A(9);
			shift_result(6) <= A(8);
			shift_result(5) <= A(7);
			shift_result(4) <= A(6);
			shift_result(3) <= A(5);
			shift_result(2) <= A(4);
			shift_result(1) <= A(3);
			shift_result(0) <= A(2);
			shifted_out <= A(1);
		end if;
		if B = "0011" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(14);
			shift_result(10) <= A(13);
			shift_result(9) <= A(12);
			shift_result(8) <= A(11);
			shift_result(7) <= A(10);
			shift_result(6) <= A(9);
			shift_result(5) <= A(8);
			shift_result(4) <= A(7);
			shift_result(3) <= A(6);
			shift_result(2) <= A(5);
			shift_result(1) <= A(4);
			shift_result(0) <= A(3);
			shifted_out <= A(2);
		end if;
		if B = "0100" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(14);
			shift_result(9) <= A(13);
			shift_result(8) <= A(12);
			shift_result(7) <= A(11);
			shift_result(6) <= A(10);
			shift_result(5) <= A(9);
			shift_result(4) <= A(8);
			shift_result(3) <= A(7);
			shift_result(2) <= A(6);
			shift_result(1) <= A(5);
			shift_result(0) <= A(4);
			shifted_out <= A(3);
		end if;
		if B = "0101" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(14);
			shift_result(8) <= A(13);
			shift_result(7) <= A(12);
			shift_result(6) <= A(11);
			shift_result(5) <= A(10);
			shift_result(4) <= A(9);
			shift_result(3) <= A(8);
			shift_result(2) <= A(7);
			shift_result(1) <= A(6);
			shift_result(0) <= A(5);
			shifted_out <= A(4);
		end if;
		if B = "0110" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(14);
			shift_result(7) <= A(13);
			shift_result(6) <= A(12);
			shift_result(5) <= A(11);
			shift_result(4) <= A(10);
			shift_result(3) <= A(9);
			shift_result(2) <= A(8);
			shift_result(1) <= A(7);
			shift_result(0) <= A(6);
			shifted_out <= A(5);
		end if;
		if B = "0111" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(14);
			shift_result(6) <= A(13);
			shift_result(5) <= A(12);
			shift_result(4) <= A(11);
			shift_result(3) <= A(10);
			shift_result(2) <= A(9);
			shift_result(1) <= A(8);
			shift_result(0) <= A(7);
			shifted_out <= A(6);
		end if;
		if B = "1000" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(14);
			shift_result(5) <= A(13);
			shift_result(4) <= A(12);
			shift_result(3) <= A(11);
			shift_result(2) <= A(10);
			shift_result(1) <= A(9);
			shift_result(0) <= A(8);
			shifted_out <= A(7);
		end if;
		if B = "1001" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(14);
			shift_result(4) <= A(13);
			shift_result(3) <= A(12);
			shift_result(2) <= A(11);
			shift_result(1) <= A(10);
			shift_result(0) <= A(9);
			shifted_out <= A(8);
		end if;
		if B = "1010" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(15);
			shift_result(4) <= A(14);
			shift_result(3) <= A(13);
			shift_result(2) <= A(12);
			shift_result(1) <= A(11);
			shift_result(0) <= A(10);
			shifted_out <= A(9);
		end if;
		if B = "1011" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(15);
			shift_result(4) <= A(15);
			shift_result(3) <= A(14);
			shift_result(2) <= A(13);
			shift_result(1) <= A(12);
			shift_result(0) <= A(11);
			shifted_out <= A(10);
		end if;
		if B = "1100" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(15);
			shift_result(4) <= A(15);
			shift_result(3) <= A(15);
			shift_result(2) <= A(14);
			shift_result(1) <= A(13);
			shift_result(0) <= A(12);
			shifted_out <= A(11);
		end if;
		if B = "1101" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(15);
			shift_result(4) <= A(15);
			shift_result(3) <= A(15);
			shift_result(2) <= A(15);
			shift_result(1) <= A(14);
			shift_result(0) <= A(13);
			shifted_out <= A(12);
		end if;
		if B = "1110" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(15);
			shift_result(4) <= A(15);
			shift_result(3) <= A(15);
			shift_result(2) <= A(15);
			shift_result(1) <= A(15);
			shift_result(0) <= A(14);
			shifted_out <= A(13);
		end if;
		if B = "1111" then
			shift_result(15) <= A(15);
			shift_result(14) <= A(15);
			shift_result(13) <= A(15);
			shift_result(12) <= A(15);
			shift_result(11) <= A(15);
			shift_result(10) <= A(15);
			shift_result(9) <= A(15);
			shift_result(8) <= A(15);
			shift_result(7) <= A(15);
			shift_result(6) <= A(15);
			shift_result(5) <= A(15);
			shift_result(4) <= A(15);
			shift_result(3) <= A(15);
			shift_result(2) <= A(15);
			shift_result(1) <= A(15);
			shift_result(0) <= A(15);
			shifted_out <= A(14);
		end if;




		else 
			shifted_out <= '0';
	end if;


	-----------------
	end process;
	
end Behavioral;
